library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;


entity rom is 
	generic (words: integer :=64;
		bits: integer :=18);
	port(
		addr: in std_logic_vector(5 downto 0);
		data: out std_logic_vector(bits-1 downto 0) );
end rom;

architecture rom_arch of rom is
	type vector_array is array(0 to words-1) of std_logic_vector(bits-1 downto 0);
	constant memory: vector_array:=(
	                --fetch 
	                "000001110000000001",
									"000110000000000010",
									"111100000000000011",
									"000010010010000000",
									
									--indirect
									"000100000000000101",
									"111100000000000110",
									"000010010011000000",
									"000000000000000000",
									--add
									"000000000101000100",
									"000100000000001010",
									"111100000000001011",
									"001000000000000000",
									--and
									"000000000101000100",
									"000100000000001110",
									"111100000000001111",
									"001100000000000000",
									--or
									"000000000101000100",
									"000100000000010010",
									"111100000000010011",
									"010000000000000000",
									--nor
									"000000000101000100",
									"000100000000010110",
									"111100000000010111",
									"010100000000000000",
									--nand
									"000000000101000100",
									"000100000000011010",
									"111100000000011011",
									"011000000000000000",
									--xor
									"000000000101000100",
									"000100000000011110",
									"111100000000011111",
									"011100000000000000",
									--xnor
									"000000000101000100",
									"000100000000100010",
									"111100000000100011",
									"100000000000000000",
									--cla
									"100100000000000000",
									"000000000000000000",
									"000000000000000000",
									"000000000000000000",
									--inca
									"000000010000000000",
									"000000000000000000",
									"000000000000000000",
									"000000000000000000",
									--sta
									"000000000101000100",
									"000000100000101110",
									"000000110000000000",
									"000000000000000000",
									--lda
									"000000000101000100",
									"000100000000110010",
									"111100000000110011",
									"000001000000000000",
									--bun
									"000000000101000100",
									"000010100000000000",
									"000000000000000000",
									"000000000000000000",
									--bsa
									"000001010000111001",
									"000000000101000100",
									"000010100000000000",
									"000000000000000000",
									--ret
									"000001100000000000",
									"000000000000000000",
									"000000000000000000",
									"000000000000000000");
	

begin
	data<=memory(conv_integer(addr));
end architecture;
